--  Analyse: ghdl -a t14_CaseWhenTb.vhdl
--  Run    : ghdl -r t14_CaseWhenTb --vcd=./t14_CaseWhenTb.vcd --stop-time=100ns
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity T14_CaseWhenTb is
end entity;

architecture behav of T14_CaseWhenTb is
    signal Sig1 : unsigned (7 downto 0) := X"AA";
    signal Sig2 : unsigned (7 downto 0) := X"BB";
    signal Sig3 : unsigned (7 downto 0) := X"CC";
    signal Sig4 : unsigned (7 downto 0) := X"DD";

    signal Sel  : unsigned (1 downto 0) := (others => '0');

    signal Output1 : unsigned (7 downto 0);
    signal Output2 : unsigned (7 downto 0);
begin
    --  Stimuli: For the sellector signal.
    process
    begin
        wait for 10 ns;
        Sel <= Sel + 1;
        wait for 10 ns;
        Sel <= Sel + 1;
        wait for 10 ns;
        Sel <= Sel + 1;
        wait for 10 ns;
        Sel <= Sel + 1;
        wait for 10 ns;
        Sel <= "UU";
        wait;
    end process;

    --  MUX using if-then-else
    process (Sel, Sig1, Sig2, Sig3, Sig4) is
    begin
        if Sel = "00" then
            Output1 <= Sig1;
        elsif Sel = "01" then
            Output1 <= Sig2;
        elsif Sel = "10" then
            Output1 <= Sig3;
        elsif Sel = "11" then
            Output1 <= Sig4;
        else --  U/X/-/etc.
            Output1 <= (others => 'X');
        end if;
    end process;


    --  MUX using case-is
    process (Sel, Sig1, Sig2, Sig3, Sig4) is
    begin
        case Sel is
            when "00" =>
                Output2 <= Sig1;

            when "01" =>
                Output2 <= Sig2;

            when "10" =>
                Output2 <= Sig3;

            when "11" =>
                Output2 <= Sig4;

            when others => --  U/X/-/etc.
                Output2 <= (others => 'X');
        end case;
    end process;
end architecture;
