--  Analyse: ghdl -a t16_GenericMux.vhdl
--  Analyse: ghdl -a t16_GenericMuxTb.vhdl
--  Run    : ghdl -r t16_GenericMuxTb --vcd=./t16_GenericMuxTb.vcd --stop-time=100ns
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity T16_GenericMuxTb is
end entity;

architecture sim of T16_GenericMuxTb is
    constant DataWidth : integer := 8;

    signal Sig1 : unsigned (DataWidth - 1 downto 0) := X"AA";
    signal Sig2 : unsigned (DataWidth - 1 downto 0) := X"BB";
    signal Sig3 : unsigned (DataWidth - 1 downto 0) := X"CC";
    signal Sig4 : unsigned (DataWidth - 1 downto 0) := X"DD";

    signal Sel  : unsigned (1 downto 0) := (others => '0');

    signal Output : unsigned (DataWidth - 1 downto 0);
begin
    --  An instance of the T16_GenericMux with architecture rtl.
    i_Mux1 : entity work.T16_GenericMux (rtl)
    generic map (
        DataWidth => DataWidth
    )
    port map (
        --  T15_Mux port => Local signal.
        Sel    => Sel,
        Sig1   => Sig1,
        Sig2   => Sig2,
        Sig3   => Sig3,
        Sig4   => Sig4,
        Output => Output
    );

    --  Testbench process.
    process
    begin
        wait for 10 ns;
        Sel <= Sel + 1;
        wait for 10 ns;
        Sel <= Sel + 1;
        wait for 10 ns;
        Sel <= Sel + 1;
        wait for 10 ns;
        Sel <= Sel + 1;
        wait for 10 ns;
        Sel <= "UU";
        wait;
    end process;
end architecture;
