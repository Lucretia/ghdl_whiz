--  Analyse: ghdl -a t09_SensitivityListTb.vhdl
--  Run    : ghdl -r t09_SensitivityListTb --stop-time=200n
entity T09_SensitivityListTb is
end entity;

architecture behav of T09_SensitivityListTb is
    signal CountUp   : Integer := 0;
    signal CountDown : Integer := 10;
begin
    process
    begin
        CountUp   <= CountUp + 1;
        CountDown <= CountDown - 1;

        wait for 10 ns;
    end process;

    --  Process triggered by "wait on"
    process
    begin
        if CountUp = CountDown then
            report "Process A: Jackpot";
        end if;

        wait on CountUp, CountDown;
    end process;

    --  Logically equivalent to A using a sensitivity list.
    process (CountUp, CountDown) is
    begin
        if CountUp = CountDown then
            report "Process B: Jackpot";
        end if;
    end process;
end architecture;
